.title KiCad schematic
R1 Net-_U1-SDA/SDI_ SDA/SDI 22
U1 __U1
R2 Net-_U1-SCL/SCK_ SCL/SCK 22
C1 +3.3V GND 100n
C2 +3.3V GND 100n
J1 __J1
D3 __D3
D4 __D4
D1 __D1
D2 __D2
.end
